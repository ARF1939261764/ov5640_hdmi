`ifndef __HDMI_CONTROLLER_CONFIG_V
`define __HDMI_CONTROLLER_CONFIG_V

/****************************************************************************************
选择FPGA型号,将通过该选项对内部的RAM进行适配
可选项：
	FPGA_TYPE_ALTERA_CYCLONE10LP
****************************************************************************************/
`define FPGA_TYPE_ALTERA_CYCLONE10LP

`endif