`ifndef __AVL_BUS_DEFINE_SV
`define __AVL_BUS_DEFINE_SV

`define ALV_BURST_MAX_COUNT           (256)

`endif
