`include "hdmi_controller_config.sv"
