module ov5640_config_data #(
  parameter DEPTH = 512
)(
  input  logic                     clk,
  input  logic[$clog2(DEPTH)-1:0]  address,
  output logic[31:0]               read_data,
  output logic[15:0]               config_data_num
);

logic[31:0] rom[DEPTH-1:0];

always @(posedge clk) begin
  read_data <= rom[address[$clog2(DEPTH)-1:0]];
end

assign rom[16'd000] = {8'h78 , 16'h3103 , 8'h11};// system clock from pad, bit[1]
assign rom[16'd001] = {8'h78 , 16'h3008 , 8'h82};// software reset, bit[7]// delay 5ms
assign rom[16'd002] = {8'h78 , 16'h3008 , 8'h42};// software power down, bit[6]
assign rom[16'd003] = {8'h78 , 16'h3103 , 8'h03};// system clock from PLL, bit[1]
assign rom[16'd004] = {8'h78 , 16'h3017 , 8'hff};// FREX, Vsync, HREF, PCLK, D[9:6] output enable
assign rom[16'd005] = {8'h78 , 16'h3018 , 8'hff};// D[5:0], GPIO[1:0] output enable
assign rom[16'd006] = {8'h78 , 16'h3034 , 8'h1A};// MIPI 10-bit
assign rom[16'd007] = {8'h78 , 16'h3037 , 8'h13};// PLL root divider, bit[4], PLL pre-divider, bit[3:0]
assign rom[16'd008] = {8'h78 , 16'h3108 , 8'h01};// PCLK root divider, bit[5:4], SCLK2x root divider, bit[3:2] // SCLK root divider, bit[1:0]
assign rom[16'd009] = {8'h78 , 16'h3630 , 8'h36};
assign rom[16'd010] = {8'h78 , 16'h3631 , 8'h0e};
assign rom[16'd011] = {8'h78 , 16'h3632 , 8'he2};
assign rom[16'd012] = {8'h78 , 16'h3633 , 8'h12};
assign rom[16'd013] = {8'h78 , 16'h3621 , 8'he0};
assign rom[16'd014] = {8'h78 , 16'h3704 , 8'ha0};
assign rom[16'd015] = {8'h78 , 16'h3703 , 8'h5a};
assign rom[16'd016] = {8'h78 , 16'h3715 , 8'h78};
assign rom[16'd017] = {8'h78 , 16'h3717 , 8'h01};
assign rom[16'd018] = {8'h78 , 16'h370b , 8'h60};
assign rom[16'd019] = {8'h78 , 16'h3705 , 8'h1a};
assign rom[16'd020] = {8'h78 , 16'h3905 , 8'h02};
assign rom[16'd021] = {8'h78 , 16'h3906 , 8'h10};
assign rom[16'd022] = {8'h78 , 16'h3901 , 8'h0a};
assign rom[16'd023] = {8'h78 , 16'h3731 , 8'h12};
assign rom[16'd024] = {8'h78 , 16'h3600 , 8'h08};// VCM control
assign rom[16'd025] = {8'h78 , 16'h3601 , 8'h33};// VCM control
assign rom[16'd026] = {8'h78 , 16'h302d , 8'h60};// system control
assign rom[16'd027] = {8'h78 , 16'h3620 , 8'h52};
assign rom[16'd028] = {8'h78 , 16'h371b , 8'h20};
assign rom[16'd029] = {8'h78 , 16'h471c , 8'h50};
assign rom[16'd030] = {8'h78 , 16'h3a13 , 8'h43};// pre-gain = 1.047x
assign rom[16'd031] = {8'h78 , 16'h3a18 , 8'h00};// gain ceiling
assign rom[16'd032] = {8'h78 , 16'h3a19 , 8'hf8};// gain ceiling = 15.5x
assign rom[16'd033] = {8'h78 , 16'h3635 , 8'h13};
assign rom[16'd034] = {8'h78 , 16'h3636 , 8'h03};
assign rom[16'd035] = {8'h78 , 16'h3634 , 8'h40};
assign rom[16'd036] = {8'h78 , 16'h3622 , 8'h01}; // 50/60Hz detection     50/60Hz 灯光条纹过滤
assign rom[16'd037] = {8'h78 , 16'h3c01 , 8'h34};// Band auto, bit[7]
assign rom[16'd038] = {8'h78 , 16'h3c04 , 8'h28};// threshold low sum
assign rom[16'd039] = {8'h78 , 16'h3c05 , 8'h98};// threshold high sum
assign rom[16'd040] = {8'h78 , 16'h3c06 , 8'h00};// light meter 1 threshold[15:8]
assign rom[16'd041] = {8'h78 , 16'h3c07 , 8'h08};// light meter 1 threshold[7:0]
assign rom[16'd042] = {8'h78 , 16'h3c08 , 8'h00};// light meter 2 threshold[15:8]
assign rom[16'd043] = {8'h78 , 16'h3c09 , 8'h1c};// light meter 2 threshold[7:0]
assign rom[16'd044] = {8'h78 , 16'h3c0a , 8'h9c};// sample number[15:8]
assign rom[16'd045] = {8'h78 , 16'h3c0b , 8'h40};// sample number[7:0]
assign rom[16'd046] = {8'h78 , 16'h3810 , 8'h00};// Timing Hoffset[11:8]
assign rom[16'd047] = {8'h78 , 16'h3811 , 8'h10};// Timing Hoffset[7:0]
assign rom[16'd048] = {8'h78 , 16'h3812 , 8'h00};// Timing Voffset[10:8]
assign rom[16'd049] = {8'h78 , 16'h3708 , 8'h64};
assign rom[16'd050] = {8'h78 , 16'h4001 , 8'h02};// BLC start from line 2
assign rom[16'd051] = {8'h78 , 16'h4005 , 8'h1a};// BLC always update
assign rom[16'd052] = {8'h78 , 16'h3000 , 8'h00};// enable blocks
assign rom[16'd053] = {8'h78 , 16'h3004 , 8'hff};// enable clocks
assign rom[16'd054] = {8'h78 , 16'h300e , 8'h58};// MIPI power down, DVP enable
assign rom[16'd055] = {8'h78 , 16'h302e , 8'h00};
assign rom[16'd056] = {8'h78 , 16'h4300 , 8'h60};// RGB565
assign rom[16'd057] = {8'h78 , 16'h501f , 8'h01};// ISP RGB
assign rom[16'd058] = {8'h78 , 16'h440e , 8'h00};
assign rom[16'd059] = {8'h78 , 16'h5000 , 8'ha7}; // Lenc on, raw gamma on, BPC on, WPC on, CIP on // AEC target    自动曝光控制
assign rom[16'd060] = {8'h78 , 16'h3a0f , 8'h30};// stable range in high
assign rom[16'd061] = {8'h78 , 16'h3a10 , 8'h28};// stable range in low
assign rom[16'd062] = {8'h78 , 16'h3a1b , 8'h30};// stable range out high
assign rom[16'd063] = {8'h78 , 16'h3a1e , 8'h26};// stable range out low
assign rom[16'd064] = {8'h78 , 16'h3a11 , 8'h60};// fast zone high
assign rom[16'd065] = {8'h78 , 16'h3a1f , 8'h14};// fast zone low// Lens correction for ?   镜头补偿
assign rom[16'd066] = {8'h78 , 16'h5800 , 8'h23};
assign rom[16'd067] = {8'h78 , 16'h5801 , 8'h14};
assign rom[16'd068] = {8'h78 , 16'h5802 , 8'h0f};
assign rom[16'd069] = {8'h78 , 16'h5803 , 8'h0f};
assign rom[16'd070] = {8'h78 , 16'h5804 , 8'h12};
assign rom[16'd071] = {8'h78 , 16'h5805 , 8'h26};
assign rom[16'd072] = {8'h78 , 16'h5806 , 8'h0c};
assign rom[16'd073] = {8'h78 , 16'h5807 , 8'h08};
assign rom[16'd074] = {8'h78 , 16'h5808 , 8'h05};
assign rom[16'd075] = {8'h78 , 16'h5809 , 8'h05};
assign rom[16'd076] = {8'h78 , 16'h580a , 8'h08};
assign rom[16'd077] = {8'h78 , 16'h580b , 8'h0d};
assign rom[16'd078] = {8'h78 , 16'h580c , 8'h08};
assign rom[16'd079] = {8'h78 , 16'h580d , 8'h03};
assign rom[16'd080] = {8'h78 , 16'h580e , 8'h00};
assign rom[16'd081] = {8'h78 , 16'h580f , 8'h00};
assign rom[16'd082] = {8'h78 , 16'h5810 , 8'h03};
assign rom[16'd083] = {8'h78 , 16'h5811 , 8'h09};
assign rom[16'd084] = {8'h78 , 16'h5812 , 8'h07};
assign rom[16'd085] = {8'h78 , 16'h5813 , 8'h03};
assign rom[16'd086] = {8'h78 , 16'h5814 , 8'h00};
assign rom[16'd087] = {8'h78 , 16'h5815 , 8'h01};
assign rom[16'd088] = {8'h78 , 16'h5816 , 8'h03};
assign rom[16'd089] = {8'h78 , 16'h5817 , 8'h08};
assign rom[16'd090] = {8'h78 , 16'h5818 , 8'h0d};
assign rom[16'd091] = {8'h78 , 16'h5819 , 8'h08};
assign rom[16'd092] = {8'h78 , 16'h581a , 8'h05};
assign rom[16'd093] = {8'h78 , 16'h581b , 8'h06};
assign rom[16'd094] = {8'h78 , 16'h581c , 8'h08};
assign rom[16'd095] = {8'h78 , 16'h581d , 8'h0e};
assign rom[16'd096] = {8'h78 , 16'h581e , 8'h29};
assign rom[16'd097] = {8'h78 , 16'h581f , 8'h17};
assign rom[16'd098] = {8'h78 , 16'h5820 , 8'h11};
assign rom[16'd099] = {8'h78 , 16'h5821 , 8'h11};
assign rom[16'd100] = {8'h78 , 16'h5822 , 8'h15};
assign rom[16'd101] = {8'h78 , 16'h5823 , 8'h28};
assign rom[16'd102] = {8'h78 , 16'h5824 , 8'h46};
assign rom[16'd103] = {8'h78 , 16'h5825 , 8'h26};
assign rom[16'd104] = {8'h78 , 16'h5826 , 8'h08};
assign rom[16'd105] = {8'h78 , 16'h5827 , 8'h26};
assign rom[16'd106] = {8'h78 , 16'h5828 , 8'h64};
assign rom[16'd107] = {8'h78 , 16'h5829 , 8'h26};
assign rom[16'd108] = {8'h78 , 16'h582a , 8'h24};
assign rom[16'd109] = {8'h78 , 16'h582b , 8'h22};
assign rom[16'd110] = {8'h78 , 16'h582c , 8'h24};
assign rom[16'd111] = {8'h78 , 16'h582d , 8'h24};
assign rom[16'd112] = {8'h78 , 16'h582e , 8'h06};
assign rom[16'd113] = {8'h78 , 16'h582f , 8'h22};
assign rom[16'd114] = {8'h78 , 16'h5830 , 8'h40};
assign rom[16'd115] = {8'h78 , 16'h5831 , 8'h42};
assign rom[16'd116] = {8'h78 , 16'h5832 , 8'h24};
assign rom[16'd117] = {8'h78 , 16'h5833 , 8'h26};
assign rom[16'd118] = {8'h78 , 16'h5834 , 8'h24};
assign rom[16'd119] = {8'h78 , 16'h5835 , 8'h22};
assign rom[16'd120] = {8'h78 , 16'h5836 , 8'h22};
assign rom[16'd121] = {8'h78 , 16'h5837 , 8'h26};
assign rom[16'd122] = {8'h78 , 16'h5838 , 8'h44};
assign rom[16'd123] = {8'h78 , 16'h5839 , 8'h24};
assign rom[16'd124] = {8'h78 , 16'h583a , 8'h26};
assign rom[16'd125] = {8'h78 , 16'h583b , 8'h28};
assign rom[16'd126] = {8'h78 , 16'h583c , 8'h42};
assign rom[16'd127] = {8'h78 , 16'h583d , 8'hce};// lenc BR offset // AWB   自动白平衡
assign rom[16'd128] = {8'h78 , 16'h5180 , 8'hff};// AWB B block
assign rom[16'd129] = {8'h78 , 16'h5181 , 8'hf2};// AWB control
assign rom[16'd130] = {8'h78 , 16'h5182 , 8'h00};// [7:4] max local counter, [3:0] max fast counter
assign rom[16'd131] = {8'h78 , 16'h5183 , 8'h14};// AWB advanced
assign rom[16'd132] = {8'h78 , 16'h5184 , 8'h25};
assign rom[16'd133] = {8'h78 , 16'h5185 , 8'h24};
assign rom[16'd134] = {8'h78 , 16'h5186 , 8'h09};
assign rom[16'd135] = {8'h78 , 16'h5187 , 8'h09};
assign rom[16'd136] = {8'h78 , 16'h5188 , 8'h09};
assign rom[16'd137] = {8'h78 , 16'h5189 , 8'h75};
assign rom[16'd138] = {8'h78 , 16'h518a , 8'h54};
assign rom[16'd139] = {8'h78 , 16'h518b , 8'he0};
assign rom[16'd140] = {8'h78 , 16'h518c , 8'hb2};
assign rom[16'd141] = {8'h78 , 16'h518d , 8'h42};
assign rom[16'd142] = {8'h78 , 16'h518e , 8'h3d};
assign rom[16'd143] = {8'h78 , 16'h518f , 8'h56};
assign rom[16'd144] = {8'h78 , 16'h5190 , 8'h46};
assign rom[16'd145] = {8'h78 , 16'h5191 , 8'hf8};// AWB top limit
assign rom[16'd146] = {8'h78 , 16'h5192 , 8'h04};// AWB bottom limit
assign rom[16'd147] = {8'h78 , 16'h5193 , 8'h70};// red limit
assign rom[16'd148] = {8'h78 , 16'h5194 , 8'hf0};// green limit
assign rom[16'd149] = {8'h78 , 16'h5195 , 8'hf0};// blue limit
assign rom[16'd150] = {8'h78 , 16'h5196 , 8'h03};// AWB control
assign rom[16'd151] = {8'h78 , 16'h5197 , 8'h01};// local limit
assign rom[16'd152] = {8'h78 , 16'h5198 , 8'h04};
assign rom[16'd153] = {8'h78 , 16'h5199 , 8'h12};
assign rom[16'd154] = {8'h78 , 16'h519a , 8'h04};
assign rom[16'd155] = {8'h78 , 16'h519b , 8'h00};
assign rom[16'd156] = {8'h78 , 16'h519c , 8'h06};
assign rom[16'd157] = {8'h78 , 16'h519d , 8'h82};
assign rom[16'd158] = {8'h78 , 16'h519e , 8'h38};// AWB control // Gamma    伽玛曲线
assign rom[16'd159] = {8'h78 , 16'h5480 , 8'h01};// Gamma bias plus on, bit[0]
assign rom[16'd160] = {8'h78 , 16'h5481 , 8'h08};
assign rom[16'd161] = {8'h78 , 16'h5482 , 8'h14};
assign rom[16'd162] = {8'h78 , 16'h5483 , 8'h28};
assign rom[16'd163] = {8'h78 , 16'h5484 , 8'h51};
assign rom[16'd164] = {8'h78 , 16'h5485 , 8'h65};
assign rom[16'd165] = {8'h78 , 16'h5486 , 8'h71};
assign rom[16'd166] = {8'h78 , 16'h5487 , 8'h7d};
assign rom[16'd167] = {8'h78 , 16'h5488 , 8'h87};
assign rom[16'd168] = {8'h78 , 16'h5489 , 8'h91};
assign rom[16'd169] = {8'h78 , 16'h548a , 8'h9a};
assign rom[16'd170] = {8'h78 , 16'h548b , 8'haa};
assign rom[16'd171] = {8'h78 , 16'h548c , 8'hb8};
assign rom[16'd172] = {8'h78 , 16'h548d , 8'hcd};
assign rom[16'd173] = {8'h78 , 16'h548e , 8'hdd};
assign rom[16'd174] = {8'h78 , 16'h548f , 8'hea};
assign rom[16'd175] = {8'h78 , 16'h5490 , 8'h1d};// color matrix   色彩矩阵
assign rom[16'd176] = {8'h78 , 16'h5381 , 8'h1e};// CMX1 for Y
assign rom[16'd177] = {8'h78 , 16'h5382 , 8'h5b};// CMX2 for Y
assign rom[16'd178] = {8'h78 , 16'h5383 , 8'h08};// CMX3 for Y
assign rom[16'd179] = {8'h78 , 16'h5384 , 8'h0a};// CMX4 for U
assign rom[16'd180] = {8'h78 , 16'h5385 , 8'h7e};// CMX5 for U
assign rom[16'd181] = {8'h78 , 16'h5386 , 8'h88};// CMX6 for U
assign rom[16'd182] = {8'h78 , 16'h5387 , 8'h7c};// CMX7 for V
assign rom[16'd183] = {8'h78 , 16'h5388 , 8'h6c};// CMX8 for V
assign rom[16'd184] = {8'h78 , 16'h5389 , 8'h10};// CMX9 for V
assign rom[16'd185] = {8'h78 , 16'h538a , 8'h01};// sign[9]
assign rom[16'd186] = {8'h78 , 16'h538b , 8'h98}; // sign[8:1] // UV adjust   UV色彩饱和度调整
assign rom[16'd187] = {8'h78 , 16'h5580 , 8'h06};// saturation on, bit[1]
assign rom[16'd188] = {8'h78 , 16'h5583 , 8'h40};
assign rom[16'd189] = {8'h78 , 16'h5584 , 8'h10};
assign rom[16'd190] = {8'h78 , 16'h5589 , 8'h10};
assign rom[16'd191] = {8'h78 , 16'h558a , 8'h00};
assign rom[16'd192] = {8'h78 , 16'h558b , 8'hf8};
assign rom[16'd193] = {8'h78 , 16'h501d , 8'h40};// enable manual offset of contrast// CIP  锐化和降噪
assign rom[16'd194] = {8'h78 , 16'h5300 , 8'h08};// CIP sharpen MT threshold 1
assign rom[16'd195] = {8'h78 , 16'h5301 , 8'h30};// CIP sharpen MT threshold 2
assign rom[16'd196] = {8'h78 , 16'h5302 , 8'h10};// CIP sharpen MT offset 1
assign rom[16'd197] = {8'h78 , 16'h5303 , 8'h00};// CIP sharpen MT offset 2
assign rom[16'd198] = {8'h78 , 16'h5304 , 8'h08};// CIP DNS threshold 1
assign rom[16'd199] = {8'h78 , 16'h5305 , 8'h30};// CIP DNS threshold 2
assign rom[16'd200] = {8'h78 , 16'h5306 , 8'h08};// CIP DNS offset 1
assign rom[16'd201] = {8'h78 , 16'h5307 , 8'h16};// CIP DNS offset 2
assign rom[16'd202] = {8'h78 , 16'h5309 , 8'h08};// CIP sharpen TH threshold 1
assign rom[16'd203] = {8'h78 , 16'h530a , 8'h30};// CIP sharpen TH threshold 2
assign rom[16'd204] = {8'h78 , 16'h530b , 8'h04};// CIP sharpen TH offset 1
assign rom[16'd205] = {8'h78 , 16'h530c , 8'h06};// CIP sharpen TH offset 2
assign rom[16'd206] = {8'h78 , 16'h5025 , 8'h00};
assign rom[16'd207] = {8'h78 , 16'h3008 , 8'h02}; // wake up from standby, bit[6]
assign rom[16'd208] = {8'h78 , 16'h3035 , 8'h11};// PLL
assign rom[16'd209] = {8'h78 , 16'h3036 , 8'h69};// PLL
assign rom[16'd210] = {8'h78 , 16'h3c07 , 8'h08};// light meter 1 threshold [7:0]
assign rom[16'd211] = {8'h78 , 16'h3820 , 8'h41};// Sensor flip off, ISP flip on
assign rom[16'd212] = {8'h78 , 16'h3821 , 8'h01};// Sensor mirror on, ISP mirror on, H binning on
assign rom[16'd213] = {8'h78 , 16'h3814 , 8'h31};// X INC
assign rom[16'd214] = {8'h78 , 16'h3815 , 8'h31};// Y INC
assign rom[16'd215] = {8'h78 , 16'h3800 , 8'h00};// HS: X address start high byte
assign rom[16'd216] = {8'h78 , 16'h3801 , 8'h00};// HS: X address start low byte
assign rom[16'd217] = {8'h78 , 16'h3802 , 8'h00};// VS: Y address start high byte
assign rom[16'd218] = {8'h78 , 16'h3803 , 8'h04};// VS: Y address start high byte
assign rom[16'd219] = {8'h78 , 16'h3804 , 8'h0a};// HW (HE)
assign rom[16'd220] = {8'h78 , 16'h3805 , 8'h3f};// HW (HE)
assign rom[16'd221] = {8'h78 , 16'h3806 , 8'h07};// VH (VE)
assign rom[16'd222] = {8'h78 , 16'h3807 , 8'h9b};// VH (VE)
assign rom[16'd223] = {8'h78 , 16'h3808 , 8'h03};// DVPHO
assign rom[16'd224] = {8'h78 , 16'h3809 , 8'h20};// DVPHO
assign rom[16'd225] = {8'h78 , 16'h380a , 8'h02};// DVPVO
assign rom[16'd226] = {8'h78 , 16'h380b , 8'h58};// DVPVO
assign rom[16'd227] = {8'h78 , 16'h380c , 8'h07};// HTS            //Total horizontal size 800
assign rom[16'd228] = {8'h78 , 16'h380d , 8'h68};// HTS
assign rom[16'd229] = {8'h78 , 16'h380e , 8'h03};// VTS            //total vertical size 500
assign rom[16'd230] = {8'h78 , 16'h380f , 8'hd8};// VTS
assign rom[16'd231] = {8'h78 , 16'h3813 , 8'h06};// Timing Voffset
assign rom[16'd232] = {8'h78 , 16'h3618 , 8'h00};
assign rom[16'd233] = {8'h78 , 16'h3612 , 8'h29};
assign rom[16'd234] = {8'h78 , 16'h3709 , 8'h52};
assign rom[16'd235] = {8'h78 , 16'h370c , 8'h03};
assign rom[16'd236] = {8'h78 , 16'h3a02 , 8'h17};// 60Hz max exposure, night mode 5fps
assign rom[16'd237] = {8'h78 , 16'h3a03 , 8'h10};// 60Hz max exposure // banding filters are calculated automatically in camera driver
assign rom[16'd238] = {8'h78 , 16'h3a14 , 8'h17};// 50Hz max exposure, night mode 5fps
assign rom[16'd239] = {8'h78 , 16'h3a15 , 8'h10};// 50Hz max exposure
assign rom[16'd240] = {8'h78 , 16'h4004 , 8'h02};// BLC 2 lines
assign rom[16'd241] = {8'h78 , 16'h3002 , 8'h1c};// reset JFIFO, SFIFO, JPEG
assign rom[16'd242] = {8'h78 , 16'h3006 , 8'hc3};// disable clock of JPEG2x, JPEG
assign rom[16'd243] = {8'h78 , 16'h4713 , 8'h03};// JPEG mode 3
assign rom[16'd244] = {8'h78 , 16'h4407 , 8'h04};// Quantization scale
assign rom[16'd245] = {8'h78 , 16'h460b , 8'h35};
assign rom[16'd246] = {8'h78 , 16'h460c , 8'h22};
assign rom[16'd247] = {8'h78 , 16'h4837 , 8'h22}; // DVP CLK divider
assign rom[16'd248] = {8'h78 , 16'h3824 , 8'h02}; // DVP CLK divider
assign rom[16'd249] = {8'h78 , 16'h5001 , 8'ha3}; // SDE on, scale on, UV average off, color matrix on, AWB on
assign rom[16'd250] = {8'h78 , 16'h3503 , 8'h00}; // AEC/AGC on
assign rom[16'd251] = {8'h78 , 16'h3035 , 8'h21};// PLL     input clock =24Mhz, PCLK =84Mhz
assign rom[16'd252] = {8'h78 , 16'h3036 , 8'h69};// PLL
assign rom[16'd253] = {8'h78 , 16'h3c07 , 8'h07}; // lightmeter 1 threshold[7:0]
assign rom[16'd254] = {8'h78 , 16'h3820 , 8'h47}; // flip
assign rom[16'd255] = {8'h78 , 16'h3821 , 8'h01}; // mirror
assign rom[16'd256] = {8'h78 , 16'h3814 , 8'h31}; // timing X inc
assign rom[16'd257] = {8'h78 , 16'h3815 , 8'h31}; // timing Y inc
assign rom[16'd258] = {8'h78 , 16'h3800 , 8'h00}; // HS
assign rom[16'd259] = {8'h78 , 16'h3801 , 8'h00}; // HS
assign rom[16'd260] = {8'h78 , 16'h3802 , 8'h00}; // VS
assign rom[16'd261] = {8'h78 , 16'h3803 , 8'h04}; // VS
assign rom[16'd262] = {8'h78 , 16'h3804 , 8'h0a}; // HW (HE)
assign rom[16'd263] = {8'h78 , 16'h3805 , 8'h3f}; // HW (HE)
assign rom[16'd264] = {8'h78 , 16'h3806 , 8'h07}; // VH (VE)
assign rom[16'd265] = {8'h78 , 16'h3807 , 8'h9f}; // VH (VE)
assign rom[16'd266] = {8'h78 , 16'h3808 , 8'h04}; // DVPHO     (1280)->1024
assign rom[16'd267] = {8'h78 , 16'h3809 , 8'h00}; // DVPHO     (1280)->1024
assign rom[16'd268] = {8'h78 , 16'h380a , 8'h03}; // DVPVO     (720)->
assign rom[16'd269] = {8'h78 , 16'h380b , 8'h00}; // DVPVO     (720)->
assign rom[16'd270] = {8'h78 , 16'h380c , 8'h07}; // HTS
assign rom[16'd271] = {8'h78 , 16'h380d , 8'h68}; // HTS
assign rom[16'd272] = {8'h78 , 16'h380e , 8'h03}; // VTS
assign rom[16'd273] = {8'h78 , 16'h380f , 8'hd8}; // VTS
assign rom[16'd274] = {8'h78 , 16'h3813 , 8'h04}; // timing V offset
assign rom[16'd275] = {8'h78 , 16'h3618 , 8'h00};
assign rom[16'd276] = {8'h78 , 16'h3612 , 8'h29};
assign rom[16'd277] = {8'h78 , 16'h3709 , 8'h52};
assign rom[16'd278] = {8'h78 , 16'h370c , 8'h03};
assign rom[16'd279] = {8'h78 , 16'h3a02 , 8'h02}; // 60Hz max exposure
assign rom[16'd280] = {8'h78 , 16'h3a03 , 8'he0}; // 60Hz max exposure
assign rom[16'd281] = {8'h78 , 16'h3a08 , 8'h00}; // B50 step
assign rom[16'd282] = {8'h78 , 16'h3a09 , 8'h6f}; // B50 step
assign rom[16'd283] = {8'h78 , 16'h3a0a , 8'h00}; // B60 step
assign rom[16'd284] = {8'h78 , 16'h3a0b , 8'h5c}; // B60 step
assign rom[16'd285] = {8'h78 , 16'h3a0e , 8'h06}; // 50Hz max band
assign rom[16'd286] = {8'h78 , 16'h3a0d , 8'h08}; // 60Hz max band
assign rom[16'd287] = {8'h78 , 16'h3a14 , 8'h02}; // 50Hz max exposure
assign rom[16'd288] = {8'h78 , 16'h3a15 , 8'he0}; // 50Hz max exposure
assign rom[16'd289] = {8'h78 , 16'h4004 , 8'h02}; // BLC line number
assign rom[16'd290] = {8'h78 , 16'h3002 , 8'h1c}; // reset JFIFO, SFIFO, JPG
assign rom[16'd291] = {8'h78 , 16'h3006 , 8'hc3}; // disable clock of JPEG2x, JPEG
assign rom[16'd292] = {8'h78 , 16'h4713 , 8'h03}; // JPEG mode 3
assign rom[16'd293] = {8'h78 , 16'h4407 , 8'h04}; // Quantization sacle
assign rom[16'd294] = {8'h78 , 16'h460b , 8'h37};
assign rom[16'd295] = {8'h78 , 16'h460c , 8'h20};
assign rom[16'd296] = {8'h78 , 16'h4837 , 8'h16}; // MIPI global timing
assign rom[16'd297] = {8'h78 , 16'h3824 , 8'h04}; // PCLK manual divider
assign rom[16'd298] = {8'h78 , 16'h3503 , 8'h00}; // AEC/AGC on
assign rom[16'd299] = {8'h78 , 16'h3016 , 8'h02}; //Strobe output enable
assign rom[16'd300] = {8'h78 , 16'h3b07 , 8'h0a}; //FREX strobe mode1
assign rom[16'd301] = {8'h78 , 16'h3b00 , 8'h83}; //STROBE CTRL: strobe request ON, Strobe mode: LED3
assign rom[16'd302] = {8'h78 , 16'h3b00 , 8'h00}; //STROBE CTRL: strobe request OFF

assign config_data_num = 303;

endmodule
