module ov5640_config(

);

endmodule
