`include "hdmi_controller_config.sv"

`define VIDEO_1024_768



